lpm_or1_inst : lpm_or1 PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		data10	 => data10_sig,
		data11	 => data11_sig,
		data12	 => data12_sig,
		data13	 => data13_sig,
		data14	 => data14_sig,
		data15	 => data15_sig,
		data16	 => data16_sig,
		data17	 => data17_sig,
		data18	 => data18_sig,
		data19	 => data19_sig,
		data2	 => data2_sig,
		data20	 => data20_sig,
		data21	 => data21_sig,
		data22	 => data22_sig,
		data23	 => data23_sig,
		data24	 => data24_sig,
		data25	 => data25_sig,
		data3	 => data3_sig,
		data4	 => data4_sig,
		data5	 => data5_sig,
		data6	 => data6_sig,
		data7	 => data7_sig,
		data8	 => data8_sig,
		data9	 => data9_sig,
		result	 => result_sig
	);
