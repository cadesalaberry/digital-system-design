lpm_or0_inst : lpm_or0 PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		result	 => result_sig
	);
