lpm_or2_inst : lpm_or2 PORT MAP (
		data0x	 => data0x_sig,
		result	 => result_sig
	);
